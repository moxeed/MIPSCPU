module programCounter(nextAddr,clk,currAddr);
input [31:0] nextAddr;
input clk;
output reg [31:0] currAddr;
	always@(posedge clk)begin
		currAddr <= nextAddr;
	end
endmodule